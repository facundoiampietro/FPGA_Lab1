library verilog;
use verilog.vl_types.all;
entity Parte_D_vlg_check_tst is
    port(
        Z1              : in     vl_logic;
        Z2              : in     vl_logic;
        Z3              : in     vl_logic;
        Z4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Parte_D_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity restador_completo_vlg_vec_tst is
end restador_completo_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Parte_D_vlg_vec_tst is
end Parte_D_vlg_vec_tst;

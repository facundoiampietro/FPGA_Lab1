library verilog;
use verilog.vl_types.all;
entity Lab_FPGA_vlg_check_tst is
    port(
        LED             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab_FPGA_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity Lab_FPGA_vlg_vec_tst is
end Lab_FPGA_vlg_vec_tst;
